-- #################################################################################################
-- # << NEORV32 - CPU Top Entity >>                                                                #
-- # ********************************************************************************************* #
-- # NEORV32 CPU:                                                                                  #
-- # * neorv32_cpu.vhd                   - CPU top entity                                          #
-- #   * neorv32_cpu_alu.vhd             - Arithmetic/logic unit                                   #
-- #     * neorv32_cpu_cp_bitmanip.vhd   - Bit-manipulation co-processor                           #
-- #     * neorv32_cpu_cp_cfu.vhd        - Custom instructions co-processor                        #
-- #     * neorv32_cpu_cp_fpu.vhd        - Single-precision FPU co-processor                       #
-- #     * neorv32_cpu_cp_muldiv.vhd     - Integer multiplier/divider co-processor                 #
-- #     * neorv32_cpu_cp_shifter.vhd    - Base ISA shifter unit                                   #
-- #   * neorv32_cpu_bus.vhd             - Load/store unit & physical memory protection            #
-- #   * neorv32_cpu_control.vhd         - CPU control and CSR system                              #
-- #     * neorv32_cpu_decompressor.vhd  - Compressed instructions decoder                         #
-- #     * neorv32_fifo.vhd              - Instruction prefetch buffer                             #
-- #   * neorv32_cpu_regfile.vhd         - Data register file                                      #
-- # * neorv32_package.vhd               - Main CPU & Processor package file                       #
-- #                                                                                               #
-- # Check out the CPU's online documentation for more information:                                #
-- #  HQ:         https://github.com/stnolting/neorv32                                             #
-- #  Data Sheet: https://stnolting.github.io/neorv32                                              #
-- #  User Guide: https://stnolting.github.io/neorv32/ug                                           #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2022, Stephan Nolting. All rights reserved.                                     #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # The NEORV32 Processor - https://github.com/stnolting/neorv32              (c) Stephan Nolting #
-- #################################################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library neorv32;
use neorv32.neorv32_package.all;

entity neorv32_cpu is
  generic (
    -- General --
    HW_THREAD_ID                 : natural; -- hardware thread id (32-bit)
    CPU_BOOT_ADDR                : std_ulogic_vector(31 downto 0); -- cpu boot address
    CPU_DEBUG_ADDR               : std_ulogic_vector(31 downto 0); -- cpu debug mode start address
    -- RISC-V CPU Extensions --
    CPU_EXTENSION_RISCV_B        : boolean; -- implement bit-manipulation extension?
    CPU_EXTENSION_RISCV_C        : boolean; -- implement compressed extension?
    CPU_EXTENSION_RISCV_E        : boolean; -- implement embedded RF extension?
    CPU_EXTENSION_RISCV_M        : boolean; -- implement mul/div extension?
    CPU_EXTENSION_RISCV_U        : boolean; -- implement user mode extension?
    CPU_EXTENSION_RISCV_Zfinx    : boolean; -- implement 32-bit floating-point extension (using INT reg!)
    CPU_EXTENSION_RISCV_Zicsr    : boolean; -- implement CSR system?
    CPU_EXTENSION_RISCV_Zicntr   : boolean; -- implement base counters?
    CPU_EXTENSION_RISCV_Zihpm    : boolean; -- implement hardware performance monitors?
    CPU_EXTENSION_RISCV_Zifencei : boolean; -- implement instruction stream sync.?
    CPU_EXTENSION_RISCV_Zmmul    : boolean; -- implement multiply-only M sub-extension?
    CPU_EXTENSION_RISCV_Zxcfu    : boolean; -- implement custom (instr.) functions unit?
    CPU_EXTENSION_RISCV_DEBUG    : boolean; -- implement CPU debug mode?
    -- Extension Options --
    FAST_MUL_EN                  : boolean; -- use DSPs for M extension's multiplier
    FAST_SHIFT_EN                : boolean; -- use barrel shifter for shift operations
    CPU_CNT_WIDTH                : natural; -- total width of CPU cycle and instret counters (0..64)
    CPU_IPB_ENTRIES              : natural; -- entries in instruction prefetch buffer, has to be a power of 2, min 2
    -- Physical Memory Protection (PMP) --
    PMP_NUM_REGIONS              : natural; -- number of regions (0..16)
    PMP_MIN_GRANULARITY          : natural; -- minimal region granularity in bytes, has to be a power of 2, min 4 bytes
    -- Hardware Performance Monitors (HPM) --
    HPM_NUM_CNTS                 : natural; -- number of implemented HPM counters (0..29)
    HPM_CNT_WIDTH                : natural  -- total size of HPM counters (0..64)
  );
  port (
    -- global control --
    clk_i         : in  std_ulogic; -- global clock, rising edge
    rstn_i        : in  std_ulogic; -- global reset, low-active, async
    sleep_o       : out std_ulogic; -- cpu is in sleep mode when set
    debug_o       : out std_ulogic; -- cpu is in debug mode when set
    priv_o        : out std_ulogic; -- current effective privilege level
    -- instruction bus interface --
    i_bus_addr_o  : out std_ulogic_vector(data_width_c-1 downto 0); -- bus access address
    i_bus_rdata_i : in  std_ulogic_vector(data_width_c-1 downto 0); -- bus read data
    i_bus_wdata_o : out std_ulogic_vector(data_width_c-1 downto 0); -- bus write data
    i_bus_ben_o   : out std_ulogic_vector(03 downto 0); -- byte enable
    i_bus_we_o    : out std_ulogic; -- write enable
    i_bus_re_o    : out std_ulogic; -- read enable
    i_bus_ack_i   : in  std_ulogic; -- bus transfer acknowledge
    i_bus_err_i   : in  std_ulogic; -- bus transfer error
    i_bus_fence_o : out std_ulogic; -- executed FENCEI operation
    -- data bus interface --
    d_bus_addr_o  : out std_ulogic_vector(data_width_c-1 downto 0); -- bus access address
    d_bus_rdata_i : in  std_ulogic_vector(data_width_c-1 downto 0); -- bus read data
    d_bus_wdata_o : out std_ulogic_vector(data_width_c-1 downto 0); -- bus write data
    d_bus_ben_o   : out std_ulogic_vector(03 downto 0); -- byte enable
    d_bus_we_o    : out std_ulogic; -- write enable
    d_bus_re_o    : out std_ulogic; -- read enable
    d_bus_ack_i   : in  std_ulogic; -- bus transfer acknowledge
    d_bus_err_i   : in  std_ulogic; -- bus transfer error
    d_bus_fence_o : out std_ulogic; -- executed FENCE operation
    -- system time input from MTIME --
    time_i        : in  std_ulogic_vector(63 downto 0); -- current system time
    -- interrupts (risc-v compliant) --
    msw_irq_i     : in  std_ulogic;-- machine software interrupt
    mext_irq_i    : in  std_ulogic;-- machine external interrupt
    mtime_irq_i   : in  std_ulogic;-- machine timer interrupt
    -- fast interrupts (custom) --
    firq_i        : in  std_ulogic_vector(15 downto 0);
    -- debug mode (halt) request --
    db_halt_req_i : in  std_ulogic
  );
end neorv32_cpu;

architecture neorv32_cpu_rtl of neorv32_cpu is

  -- local signals --
  signal ctrl        : std_ulogic_vector(ctrl_width_c-1 downto 0); -- main control bus
  signal comparator  : std_ulogic_vector(1 downto 0); -- comparator result
  signal imm         : std_ulogic_vector(data_width_c-1 downto 0); -- immediate
  signal rs1, rs2    : std_ulogic_vector(data_width_c-1 downto 0); -- source registers
  signal alu_res     : std_ulogic_vector(data_width_c-1 downto 0); -- alu result
  signal alu_add     : std_ulogic_vector(data_width_c-1 downto 0); -- alu address result
  signal mem_rdata   : std_ulogic_vector(data_width_c-1 downto 0); -- memory read data
  signal alu_idone   : std_ulogic; -- iterative alu operation done
  signal bus_d_wait  : std_ulogic; -- wait for current bus data access
  signal csr_rdata   : std_ulogic_vector(data_width_c-1 downto 0); -- csr read data
  signal mar         : std_ulogic_vector(data_width_c-1 downto 0); -- current memory address register
  signal ma_load     : std_ulogic; -- misaligned load data address
  signal ma_store    : std_ulogic; -- misaligned store data address
  signal be_load     : std_ulogic; -- bus error on load data access
  signal be_store    : std_ulogic; -- bus error on store data access
  signal fetch_pc    : std_ulogic_vector(data_width_c-1 downto 0); -- pc for instruction fetch
  signal curr_pc     : std_ulogic_vector(data_width_c-1 downto 0); -- current pc (for current executed instruction)
  signal next_pc     : std_ulogic_vector(data_width_c-1 downto 0); -- next pc (for next executed instruction)
  signal fpu_flags   : std_ulogic_vector(4 downto 0); -- FPU exception flags
  signal i_pmp_fault : std_ulogic; -- instruction fetch PMP fault

  -- pmp interface --
  signal pmp_addr : pmp_addr_if_t;
  signal pmp_ctrl : pmp_ctrl_if_t;

begin

  -- CPU ISA Configuration ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  assert false report
  "NEORV32 CPU ISA Configuration (MARCH): " &
  cond_sel_string_f(CPU_EXTENSION_RISCV_E, "RV32E", "RV32I") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_M, "M", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_C, "C", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_B, "B", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_U, "U", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_Zicsr, "_Zicsr", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_Zicntr, "_Zicntr", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_Zihpm, "_Zihpm", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_Zifencei, "_Zifencei", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_Zfinx, "_Zfinx", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_Zmmul, "_Zmmul", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_Zxcfu, "_Zxcfu", "") &
  cond_sel_string_f(CPU_EXTENSION_RISCV_DEBUG, "_DebugMode", "") &
  ""
  severity note;


  -- Sanity Checks --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- simulation notifier --
  assert not (is_simulation_c = true)  report "NEORV32 CPU INFO: Seems like this is a simulation." severity note;
  assert not (is_simulation_c = false) report "NEORV32 CPU INFO: Seems like this is real hardware." severity note;

  -- hardware reset notifier --
  assert not (dedicated_reset_c = false) report "NEORV32 CPU CONFIG NOTE: Implementing NO dedicated hardware reset for uncritical registers (default)." severity note;
  assert not (dedicated_reset_c = true)  report "NEORV32 CPU CONFIG NOTE: Implementing defined hardware reset for uncritical registers (non-default, reset-to-zero, might increase area)." severity note;
  assert not ((def_rst_val_c /= '-') and (def_rst_val_c /= '0')) report "NEORV32 CPU CONFIG ERROR! Invalid configuration of package <def_rst_val_c> constant (has to be '-' or '0')." severity error;

  -- CPU boot address alignment --
  assert not (CPU_BOOT_ADDR(1 downto 0) /= "00") report "NEORV32 CPU CONFIG ERROR! <CPU_BOOT_ADDR> has to be 32-bit aligned." severity error;

  -- CSR system --
  assert not (CPU_EXTENSION_RISCV_Zicsr = false) report "NEORV32 CPU CONFIG WARNING! No exception/interrupt/trap/privileged features available when <CPU_EXTENSION_RISCV_Zicsr> = false." severity warning;

  -- CPU counters (cycle and instret) --
  assert not ((CPU_EXTENSION_RISCV_Zicntr = true) and ((CPU_CNT_WIDTH < 0) or (CPU_CNT_WIDTH > 64))) report "NEORV32 CPU CONFIG ERROR! Invalid <CPU_CNT_WIDTH> configuration. Has to be 0..64." severity error;
  assert not ((CPU_EXTENSION_RISCV_Zicntr = true) and (CPU_CNT_WIDTH < 64)) report "NEORV32 CPU CONFIG WARNING! Implementing CPU <cycle> and <instret> CSRs with reduced size (" & integer'image(CPU_CNT_WIDTH) & "-bit instead of 64-bit). This is not RISC-V compliant and might have unintended SW side effects." severity warning;

  -- U-extension requires Zicsr extension --
  assert not ((CPU_EXTENSION_RISCV_Zicsr = false) and (CPU_EXTENSION_RISCV_U = true)) report "NEORV32 CPU CONFIG ERROR! User mode requires <CPU_EXTENSION_RISCV_Zicsr> extension to be enabled." severity error;

  -- Instruction prefetch buffer --
  assert not (is_power_of_two_f(CPU_IPB_ENTRIES) = false) report "NEORV32 CPU CONFIG ERROR! Number of entries in instruction prefetch buffer <CPU_IPB_ENTRIES> has to be a power of two." severity error;
  assert not (CPU_IPB_ENTRIES < 2) report "NEORV32 CPU CONFIG ERROR! Number of entries in instruction prefetch buffer <CPU_IPB_ENTRIES> has to be >= 2." severity error;

  -- PMP check --
  assert not (PMP_NUM_REGIONS > 16) report "NEORV32 CPU CONFIG ERROR! Number of PMP regions <PMP_NUM_REGIONS> out of valid range (0..16)." severity error;
  assert not ((is_power_of_two_f(PMP_MIN_GRANULARITY) = false) and (PMP_NUM_REGIONS > 0)) report "NEORV32 CPU CONFIG ERROR! <PMP_MIN_GRANULARITY> has to be a power of two." severity error;
  assert not ((PMP_MIN_GRANULARITY < 4) and (PMP_NUM_REGIONS > 0)) report "NEORV32 CPU CONFIG ERROR! <PMP_MIN_GRANULARITY> has to be >= 4 bytes." severity error;
  assert not ((CPU_EXTENSION_RISCV_Zicsr = false) and (PMP_NUM_REGIONS > 0)) report "NEORV32 CPU CONFIG ERROR! Physical memory protection (PMP) requires <CPU_EXTENSION_RISCV_Zicsr> extension to be enabled." severity error;

  -- HPM counters check --
  assert not ((CPU_EXTENSION_RISCV_Zihpm = true) and (HPM_NUM_CNTS > 29)) report "NEORV32 CPU CONFIG ERROR! Number of HPM counters <HPM_NUM_CNTS> out of valid range (0..29)." severity error;
  assert not ((CPU_EXTENSION_RISCV_Zihpm = true) and ((HPM_CNT_WIDTH < 0) or (HPM_CNT_WIDTH > 64))) report "NEORV32 CPU CONFIG ERROR! HPM counter width <HPM_CNT_WIDTH> has to be 0..64 bit." severity error; 
  assert not ((CPU_EXTENSION_RISCV_Zicsr = false) and (CPU_EXTENSION_RISCV_Zihpm = true)) report "NEORV32 CPU CONFIG ERROR! Hardware performance monitors extension <CPU_EXTENSION_RISCV_Zihpm> requires <CPU_EXTENSION_RISCV_Zicsr> extension to be enabled." severity error;

  -- Mul-extension --
  assert not ((CPU_EXTENSION_RISCV_Zmmul = true) and (CPU_EXTENSION_RISCV_M = true)) report "NEORV32 CPU CONFIG ERROR! <M> and <Zmmul> extensions cannot co-exist!" severity error;

  -- Custom Functions Unit --
  assert not (CPU_EXTENSION_RISCV_Zxcfu = true) report "NEORV32 CPU CONFIG NOTE: Implementing Custom Functions Unit (CFU) as <Zxcfu> ISA extension." severity note;

  -- Debug mode --
  assert not ((CPU_EXTENSION_RISCV_DEBUG = true) and (CPU_EXTENSION_RISCV_Zicsr = false)) report "NEORV32 CPU CONFIG ERROR! Debug mode requires <CPU_EXTENSION_RISCV_Zicsr> extension to be enabled." severity error;
  assert not ((CPU_EXTENSION_RISCV_DEBUG = true) and (CPU_EXTENSION_RISCV_Zifencei = false)) report "NEORV32 CPU CONFIG ERROR! Debug mode requires <CPU_EXTENSION_RISCV_Zifencei> extension to be enabled." severity error;

  -- fast multiplication option --
  assert not (FAST_MUL_EN = true) report "NEORV32 CPU CONFIG NOTE: <FAST_MUL_EN> set. Trying to use DSP blocks for base ISA multiplications." severity note;

  -- fast shift option --
  assert not (FAST_SHIFT_EN = true) report "NEORV32 CPU CONFIG NOTE: <FAST_SHIFT_EN> set. Implementing full-parallel logic / barrel shifters." severity note;


  -- Control Unit ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  neorv32_cpu_control_inst: neorv32_cpu_control
  generic map (
    -- General --
    HW_THREAD_ID                 => HW_THREAD_ID,                 -- hardware thread id
    CPU_BOOT_ADDR                => CPU_BOOT_ADDR,                -- cpu boot address
    CPU_DEBUG_ADDR               => CPU_DEBUG_ADDR,               -- cpu debug mode start address
    -- RISC-V CPU Extensions --
    CPU_EXTENSION_RISCV_B        => CPU_EXTENSION_RISCV_B,        -- implement bit-manipulation extension?
    CPU_EXTENSION_RISCV_C        => CPU_EXTENSION_RISCV_C,        -- implement compressed extension?
    CPU_EXTENSION_RISCV_E        => CPU_EXTENSION_RISCV_E,        -- implement embedded RF extension?
    CPU_EXTENSION_RISCV_M        => CPU_EXTENSION_RISCV_M,        -- implement mul/div extension?
    CPU_EXTENSION_RISCV_U        => CPU_EXTENSION_RISCV_U,        -- implement user mode extension?
    CPU_EXTENSION_RISCV_Zfinx    => CPU_EXTENSION_RISCV_Zfinx,    -- implement 32-bit floating-point extension (using INT reg!)
    CPU_EXTENSION_RISCV_Zicsr    => CPU_EXTENSION_RISCV_Zicsr,    -- implement CSR system?
    CPU_EXTENSION_RISCV_Zicntr   => CPU_EXTENSION_RISCV_Zicntr,   -- implement base counters?
    CPU_EXTENSION_RISCV_Zihpm    => CPU_EXTENSION_RISCV_Zihpm,    -- implement hardware performance monitors?
    CPU_EXTENSION_RISCV_Zifencei => CPU_EXTENSION_RISCV_Zifencei, -- implement instruction stream sync.?
    CPU_EXTENSION_RISCV_Zmmul    => CPU_EXTENSION_RISCV_Zmmul,    -- implement multiply-only M sub-extension?
    CPU_EXTENSION_RISCV_Zxcfu    => CPU_EXTENSION_RISCV_Zxcfu,    -- implement custom (instr.) functions unit?
    CPU_EXTENSION_RISCV_DEBUG    => CPU_EXTENSION_RISCV_DEBUG,    -- implement CPU debug mode?
    -- Tuning Options --
    FAST_MUL_EN                  => FAST_MUL_EN,                  -- use DSPs for M extension's multiplier
    FAST_SHIFT_EN                => FAST_SHIFT_EN,                -- use barrel shifter for shift operations
    CPU_CNT_WIDTH                => CPU_CNT_WIDTH,                -- total width of CPU cycle and instret counters (0..64)
    CPU_IPB_ENTRIES              => CPU_IPB_ENTRIES,              -- entries is instruction prefetch buffer, has to be a power of 2, min 2
    -- Physical memory protection (PMP) --
    PMP_NUM_REGIONS              => PMP_NUM_REGIONS,              -- number of regions (0..16)
    PMP_MIN_GRANULARITY          => PMP_MIN_GRANULARITY,          -- minimal region granularity in bytes, has to be a power of 2, min 4 bytes
    -- Hardware Performance Monitors (HPM) --
    HPM_NUM_CNTS                 => HPM_NUM_CNTS,                 -- number of implemented HPM counters (0..29)
    HPM_CNT_WIDTH                => HPM_CNT_WIDTH                 -- total size of HPM counters
  )
  port map (
    -- global control --
    clk_i         => clk_i,         -- global clock, rising edge
    rstn_i        => rstn_i,        -- global reset, low-active, async
    ctrl_o        => ctrl,          -- main control bus
    -- instruction fetch interface --
    i_bus_addr_o  => fetch_pc,      -- bus access address
    i_bus_rdata_i => i_bus_rdata_i, -- bus read data
    i_bus_re_o    => i_bus_re_o,    -- read enable
    i_bus_ack_i   => i_bus_ack_i,   -- bus transfer acknowledge
    i_bus_err_i   => i_bus_err_i,   -- bus transfer error
    i_pmp_fault_i => i_pmp_fault,   -- instruction fetch pmp fault
    -- status input --
    alu_idone_i   => alu_idone,     -- ALU iterative operation done
    bus_d_wait_i  => bus_d_wait,    -- wait for bus
    -- data input --
    cmp_i         => comparator,    -- comparator status
    alu_add_i     => alu_add,       -- ALU address result
    rs1_i         => rs1,           -- rf source 1
    -- data output --
    imm_o         => imm,           -- immediate
    curr_pc_o     => curr_pc,       -- current PC (corresponding to current instruction)
    next_pc_o     => next_pc,       -- next PC (corresponding to next instruction)
    csr_rdata_o   => csr_rdata,     -- CSR read data
    -- FPU interface --
    fpu_flags_i   => fpu_flags,     -- exception flags
    -- debug mode (halt) request --
    db_halt_req_i => db_halt_req_i,
    -- interrupts (risc-v compliant) --
    msw_irq_i     => msw_irq_i,     -- machine software interrupt
    mext_irq_i    => mext_irq_i,    -- machine external interrupt
    mtime_irq_i   => mtime_irq_i,   -- machine timer interrupt
    -- fast interrupts (custom) --
    firq_i        => firq_i,        -- fast interrupt trigger
    -- system time input from MTIME --
    time_i        => time_i,        -- current system time
    -- physical memory protection --
    pmp_addr_o    => pmp_addr,      -- addresses
    pmp_ctrl_o    => pmp_ctrl,      -- configs
    -- bus access exceptions --
    mar_i         => mar,           -- memory address register
    ma_load_i     => ma_load,       -- misaligned load data address
    ma_store_i    => ma_store,      -- misaligned store data address
    be_load_i     => be_load,       -- bus error on load data access
    be_store_i    => be_store       -- bus error on store data access
  );

  -- CPU state --
  sleep_o <= ctrl(ctrl_sleep_c); -- set when CPU is sleeping (after WFI)
  debug_o <= ctrl(ctrl_debug_running_c); -- set when CPU is in debug mode
  priv_o  <= ctrl(ctrl_priv_mode_c); -- current effective privilege level

  -- instruction fetch interface --
  i_bus_addr_o  <= fetch_pc;
  i_bus_wdata_o <= (others => '0'); -- read-only
  i_bus_ben_o   <= (others => '0'); -- read-only
  i_bus_we_o    <= '0'; -- read-only
  i_bus_fence_o <= ctrl(ctrl_bus_fencei_c);


  -- Register File --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  neorv32_cpu_regfile_inst: neorv32_cpu_regfile
  generic map (
    CPU_EXTENSION_RISCV_E => CPU_EXTENSION_RISCV_E -- implement embedded RF extension?
  )
  port map (
    -- global control --
    clk_i  => clk_i,     -- global clock, rising edge
    ctrl_i => ctrl,      -- main control bus
    -- data input --
    alu_i  => alu_res,   -- ALU result
    mem_i  => mem_rdata, -- memory read data
    csr_i  => csr_rdata, -- CSR read data
    pc2_i  => next_pc,   -- next PC
    -- data output --
    rs1_o  => rs1,       -- operand 1
    rs2_o  => rs2        -- operand 2
  );


  -- ALU ------------------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  neorv32_cpu_alu_inst: neorv32_cpu_alu
  generic map (
    -- RISC-V CPU Extensions --
    CPU_EXTENSION_RISCV_B     => CPU_EXTENSION_RISCV_B,     -- implement bit-manipulation extension?
    CPU_EXTENSION_RISCV_M     => CPU_EXTENSION_RISCV_M,     -- implement mul/div extension?
    CPU_EXTENSION_RISCV_Zmmul => CPU_EXTENSION_RISCV_Zmmul, -- implement multiply-only M sub-extension?
    CPU_EXTENSION_RISCV_Zfinx => CPU_EXTENSION_RISCV_Zfinx, -- implement 32-bit floating-point extension (using INT reg!)
    CPU_EXTENSION_RISCV_Zxcfu => CPU_EXTENSION_RISCV_Zxcfu, -- implement custom (instr.) functions unit?
    -- Extension Options --
    FAST_MUL_EN               => FAST_MUL_EN,               -- use DSPs for M extension's multiplier
    FAST_SHIFT_EN             => FAST_SHIFT_EN              -- use barrel shifter for shift operations
  )
  port map (
    -- global control --
    clk_i       => clk_i,      -- global clock, rising edge
    rstn_i      => rstn_i,     -- global reset, low-active, async
    ctrl_i      => ctrl,       -- main control bus
    -- data input --
    rs1_i       => rs1,        -- rf source 1
    rs2_i       => rs2,        -- rf source 2
    pc_i        => curr_pc,    -- current PC
    imm_i       => imm,        -- immediate
    -- data output --
    cmp_o       => comparator, -- comparator status
    res_o       => alu_res,    -- ALU result
    add_o       => alu_add,    -- address computation result
    fpu_flags_o => fpu_flags,  -- FPU exception flags
    -- status --
    idone_o     => alu_idone   -- iterative processing units done?
  );


  -- Bus Interface (Load/Store Unit) --------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  neorv32_cpu_bus_inst: neorv32_cpu_bus
  generic map (
    PMP_NUM_REGIONS     => PMP_NUM_REGIONS,    -- number of regions (0..16)
    PMP_MIN_GRANULARITY => PMP_MIN_GRANULARITY -- minimal region granularity in bytes, has to be a power of 2, min 4 bytes
  )
  port map (
    -- global control --
    clk_i         => clk_i,         -- global clock, rising edge
    rstn_i        => rstn_i,        -- global reset, low-active, async
    ctrl_i        => ctrl,          -- main control bus
    -- cpu instruction fetch interface --
    fetch_pc_i    => fetch_pc,      -- PC for instruction fetch
    i_pmp_fault_o => i_pmp_fault,   -- instruction fetch pmp fault
    -- cpu data access interface --
    addr_i        => alu_add,       -- ALU.add result -> access address
    wdata_i       => rs2,           -- write data
    rdata_o       => mem_rdata,     -- read data
    mar_o         => mar,           -- current memory address register
    d_wait_o      => bus_d_wait,    -- wait for access to complete
    ma_load_o     => ma_load,       -- misaligned load data address
    ma_store_o    => ma_store,      -- misaligned store data address
    be_load_o     => be_load,       -- bus error on load data access
    be_store_o    => be_store,      -- bus error on store data access
    -- physical memory protection --
    pmp_addr_i    => pmp_addr,      -- addresses
    pmp_ctrl_i    => pmp_ctrl,      -- configurations
    -- data bus --
    d_bus_addr_o  => d_bus_addr_o,  -- bus access address
    d_bus_rdata_i => d_bus_rdata_i, -- bus read data
    d_bus_wdata_o => d_bus_wdata_o, -- bus write data
    d_bus_ben_o   => d_bus_ben_o,   -- byte enable
    d_bus_we_o    => d_bus_we_o,    -- write enable
    d_bus_re_o    => d_bus_re_o,    -- read enable
    d_bus_ack_i   => d_bus_ack_i,   -- bus transfer acknowledge
    d_bus_err_i   => d_bus_err_i,   -- bus transfer error
    d_bus_fence_o => d_bus_fence_o  -- fence operation
  );


end neorv32_cpu_rtl;
