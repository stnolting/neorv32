library ieee;
use ieee.std_logic_1164.all;

package neorv32_bootrom_image is

type rom_t is array (0 to 1023) of std_ulogic_vector(31 downto 0);
constant image_size_c : natural := 3848;
constant image_data_c : rom_t := (
x"f14020f3",
x"80200217",
x"0fb20213",
x"ff027113",
x"80200197",
x"7f018193",
x"000022b7",
x"80028293",
x"30029073",
x"00000317",
x"0ec30313",
x"30531073",
x"30401073",
x"00001397",
x"ed438393",
x"80200417",
x"fc440413",
x"80200497",
x"fbc48493",
x"80200517",
x"fb450513",
x"80200597",
x"fb458593",
x"00000613",
x"00000693",
x"00000713",
x"00000793",
x"04008263",
x"00000797",
x"01c78793",
x"30579073",
x"30445073",
x"30046073",
x"10500073",
x"ffdff06f",
x"00000797",
x"08478793",
x"30579073",
x"fff44737",
x"00872103",
x"00c72603",
x"fff40737",
x"00072223",
x"0380006f",
x"00838e63",
x"00945c63",
x"0003a783",
x"00f42023",
x"00438393",
x"00440413",
x"fedff06f",
x"00b55863",
x"00052023",
x"00450513",
x"ff5ff06f",
x"00000617",
x"73460613",
x"0ff0000f",
x"0000100f",
x"00000513",
x"00000593",
x"000600e7",
x"30047073",
x"30401073",
x"00000597",
x"01058593",
x"30559073",
x"34051073",
x"10500073",
x"ffdff06f",
x"00000513",
x"00008067",
x"fffe07b7",
x"0087a783",
x"00000513",
x"00e79713",
x"00075e63",
x"fff507b7",
x"0007a703",
x"00f71693",
x"fe06dce3",
x"0047a503",
x"0ff57513",
x"00008067",
x"ff010113",
x"00812423",
x"00912223",
x"00112623",
x"00050493",
x"00000413",
x"fb9ff0ef",
x"00440793",
x"002787b3",
x"fea78e23",
x"00140413",
x"00400793",
x"fef414e3",
x"00012783",
x"00c12083",
x"00812403",
x"00f4a023",
x"00000513",
x"00412483",
x"01010113",
x"00008067",
x"fffe07b7",
x"0087a783",
x"00e79713",
x"02075c63",
x"00a00793",
x"00f51e63",
x"fff507b7",
x"0007a703",
x"00c71693",
x"fe06dce3",
x"00d00713",
x"00e7a223",
x"fff507b7",
x"0007a703",
x"00c71693",
x"fe06dce3",
x"00a7a223",
x"00008067",
x"ff810113",
x"00812023",
x"00112223",
x"00050413",
x"00044503",
x"00051a63",
x"00412083",
x"00012403",
x"00810113",
x"00008067",
x"00140413",
x"f8dff0ef",
x"fe1ff06f",
x"fdc10113",
x"00812e23",
x"00912c23",
x"02112023",
x"800004b7",
x"00058413",
x"0004a223",
x"000500e7",
x"02050663",
x"ffe01537",
x"c8450513",
x"fa1ff0ef",
x"00100793",
x"02012083",
x"01c12403",
x"01812483",
x"00078513",
x"02410113",
x"00008067",
x"01410513",
x"00012a23",
x"00012823",
x"00012623",
x"000400e7",
x"00a12023",
x"01010513",
x"000400e7",
x"00a12223",
x"00c10513",
x"000400e7",
x"01412703",
x"b007c7b7",
x"0de78793",
x"00f70863",
x"ffe01537",
x"c9850513",
x"f9dff06f",
x"00412703",
x"00012783",
x"00012423",
x"00e7e7b3",
x"00a7e7b3",
x"00000713",
x"01012683",
x"02d77c63",
x"f60798e3",
x"00810513",
x"00e12023",
x"000400e7",
x"00c12683",
x"00812603",
x"00012703",
x"00050793",
x"00c686b3",
x"00d12623",
x"00c72023",
x"00470713",
x"fc9ff06f",
x"f2079ee3",
x"00c12603",
x"fff00713",
x"00e60863",
x"ffe01537",
x"cac50513",
x"f2dff06f",
x"ffe01537",
x"cc050513",
x"00f12023",
x"00d4a223",
x"eb9ff0ef",
x"0ff0000f",
x"00012783",
x"f15ff06f",
x"ff410113",
x"00912023",
x"00050493",
x"03000513",
x"00112423",
x"00812223",
x"e49ff0ef",
x"07800513",
x"e41ff0ef",
x"01c00413",
x"0084d733",
x"ffe017b7",
x"00f77713",
x"ef878793",
x"00e787b3",
x"0007c503",
x"ffc40413",
x"e1dff0ef",
x"ffc00793",
x"fcf41ee3",
x"00812083",
x"00412403",
x"00012483",
x"00c10113",
x"00008067",
x"fff4c7b7",
x"ffc7a583",
x"ff87a503",
x"ffc7a703",
x"fee59ae3",
x"00008067",
x"fff80737",
x"00072783",
x"00d79693",
x"fe06cce3",
x"800007b7",
x"00878793",
x"00f72223",
x"00008067",
x"fff807b7",
x"0007a703",
x"00d71693",
x"fe06cce3",
x"80000737",
x"00e7a223",
x"00008067",
x"fff807b7",
x"00a7a223",
x"0007a703",
x"fe074ee3",
x"0047a503",
x"0ff57513",
x"00008067",
x"ff810113",
x"00112223",
x"00a12023",
x"f9dff0ef",
x"00012503",
x"fd1ff0ef",
x"00412083",
x"00810113",
x"fa9ff06f",
x"ff810113",
x"00112223",
x"f7dff0ef",
x"00500513",
x"fb1ff0ef",
x"00000513",
x"fa9ff0ef",
x"00a12023",
x"f85ff0ef",
x"00412083",
x"00012503",
x"00810113",
x"00008067",
x"fffe07b7",
x"0087a783",
x"00100513",
x"00d79713",
x"06075463",
x"ffc10113",
x"00112023",
x"fff807b7",
x"0007a023",
x"01900713",
x"00e7a023",
x"0ab00513",
x"800007b7",
x"00400737",
x"00e7a023",
x"f6dff0ef",
x"00600513",
x"f65ff0ef",
x"f85ff0ef",
x"00257793",
x"fff00513",
x"00078c63",
x"00400513",
x"f4dff0ef",
x"f6dff0ef",
x"01e51793",
x"41f7d513",
x"00012083",
x"00410113",
x"00008067",
x"00008067",
x"ff810113",
x"800007b7",
x"00812023",
x"0007a403",
x"00112223",
x"01045513",
x"0ff57513",
x"ef5ff0ef",
x"00845513",
x"0ff57513",
x"ee9ff0ef",
x"0ff47513",
x"00012403",
x"00412083",
x"00810113",
x"ed5ff06f",
x"ff010113",
x"00112623",
x"00812423",
x"00912223",
x"00050493",
x"e81ff0ef",
x"00300513",
x"eb5ff0ef",
x"fa1ff0ef",
x"00000413",
x"00000513",
x"ea5ff0ef",
x"00440793",
x"002787b3",
x"fea78e23",
x"00140413",
x"00400793",
x"fef412e3",
x"e6dff0ef",
x"00012783",
x"80000737",
x"00c12083",
x"00f4a023",
x"00072783",
x"00412483",
x"00000513",
x"008787b3",
x"00812403",
x"00f72023",
x"01010113",
x"00008067",
x"ff410113",
x"00812223",
x"00112423",
x"00a12023",
x"00000413",
x"00600513",
x"e59ff0ef",
x"dfdff0ef",
x"00200513",
x"e31ff0ef",
x"f1dff0ef",
x"00440793",
x"002787b3",
x"ffc7c503",
x"e1dff0ef",
x"dfdff0ef",
x"e55ff0ef",
x"00157513",
x"fe051ce3",
x"80000737",
x"00072783",
x"00140413",
x"00178793",
x"00f72023",
x"00400793",
x"faf418e3",
x"00812083",
x"00412403",
x"00c10113",
x"00008067",
x"fd410113",
x"02112423",
x"02512223",
x"02612023",
x"00712e23",
x"00812c23",
x"00a12a23",
x"00b12823",
x"00c12623",
x"00d12423",
x"00e12223",
x"00f12023",
x"34202473",
x"800007b7",
x"00778793",
x"fffe0737",
x"08f41e63",
x"00872783",
x"01079713",
x"00075a63",
x"fffc0737",
x"00472783",
x"0017c793",
x"00f72223",
x"fffe0437",
x"00842783",
x"00f79713",
x"02075e63",
x"d19ff0ef",
x"00042783",
x"0027d793",
x"00a78533",
x"00f537b3",
x"00b787b3",
x"f1402773",
x"fff446b7",
x"00371713",
x"00d70733",
x"fff00693",
x"00d72023",
x"00f72223",
x"00a72023",
x"01812403",
x"02812083",
x"02412283",
x"02012303",
x"01c12383",
x"01412503",
x"01012583",
x"00c12603",
x"00812683",
x"00412703",
x"00012783",
x"02c10113",
x"30200073",
x"00872783",
x"00e79713",
x"04075a63",
x"ffe01537",
x"cc450513",
x"addff0ef",
x"00040513",
x"c2dff0ef",
x"02000513",
x"a85ff0ef",
x"34102573",
x"c1dff0ef",
x"02000513",
x"a75ff0ef",
x"34a02573",
x"c0dff0ef",
x"02000513",
x"a65ff0ef",
x"34302573",
x"bfdff0ef",
x"ffe01537",
x"ce050513",
x"a99ff0ef",
x"fffe07b7",
x"0087a783",
x"01079713",
x"00075863",
x"fffc07b7",
x"00100713",
x"00e7a223",
x"99dff06f",
x"800007b7",
x"0047a783",
x"ffc10113",
x"00112023",
x"00079e63",
x"ffe01537",
x"ce850513",
x"a59ff0ef",
x"989ff0ef",
x"07900793",
x"06f51263",
x"000027b7",
x"80078793",
x"30079073",
x"fffe07b7",
x"0087a783",
x"01079713",
x"00075663",
x"fffc07b7",
x"0007a223",
x"ffe01537",
x"d0c50513",
x"a1dff0ef",
x"00000513",
x"b6dff0ef",
x"ffe01537",
x"d1c50513",
x"a09ff0ef",
x"fff50737",
x"00072783",
x"fe07cee3",
x"00000793",
x"0000100f",
x"34179073",
x"30200073",
x"00012083",
x"00410113",
x"00008067",
x"fec10113",
x"ffe007b7",
x"00112823",
x"00812623",
x"00912423",
x"62078793",
x"30579073",
x"fffe07b7",
x"0087a703",
x"01071693",
x"0006d863",
x"fffc0737",
x"00100693",
x"00d72223",
x"0087a703",
x"00e71693",
x"0406dc63",
x"fff50737",
x"00072023",
x"ffff7637",
x"00009737",
x"0007a683",
x"5ff70713",
x"00000793",
x"a0060613",
x"12d76663",
x"00000713",
x"3fe00613",
x"12f66663",
x"fff78793",
x"3ff7f793",
x"00371713",
x"01877713",
x"00679793",
x"00e7e7b3",
x"0017e793",
x"fff50737",
x"00f72023",
x"fffe07b7",
x"0087a703",
x"00f71693",
x"0206da63",
x"fff4c737",
x"fe072c23",
x"fe072e23",
x"0007a783",
x"fff44737",
x"0027d793",
x"00f72023",
x"00072223",
x"08000793",
x"30479073",
x"00800793",
x"3007a073",
x"ffe01537",
x"d2450513",
x"8fdff0ef",
x"ffe01537",
x"d5050513",
x"8f1ff0ef",
x"fffe0437",
x"00842783",
x"00f79713",
x"0c075863",
x"ffe01537",
x"d5c50513",
x"8d5ff0ef",
x"a8dff0ef",
x"00042403",
x"00341413",
x"00a404b3",
x"0084b433",
x"00b40433",
x"fffe07b7",
x"0087a783",
x"00e79713",
x"08075663",
x"fff507b7",
x"0007a703",
x"00f71693",
x"0606de63",
x"ffe01537",
x"0047a783",
x"d8050513",
x"88dff0ef",
x"ffe01537",
x"db450513",
x"881ff0ef",
x"ffe01537",
x"dc850513",
x"875ff0ef",
x"fa4ff0ef",
x"00050413",
x"821ff0ef",
x"00a00513",
x"819ff0ef",
x"07200793",
x"06f41e63",
x"ffe002b7",
x"00028067",
x"00c686b3",
x"00178793",
x"ecdff06f",
x"ffe70693",
x"ffd6f693",
x"00069863",
x"0037d793",
x"00170713",
x"ec1ff06f",
x"0017d793",
x"ff5ff06f",
x"9ddff0ef",
x"f685e2e3",
x"00b41463",
x"f4956ee3",
x"00a00513",
x"fc4ff0ef",
x"ffe01537",
x"d8c50513",
x"801ff0ef",
x"ffe005b7",
x"ffe00537",
x"52c58593",
x"47050513",
x"821ff0ef",
x"f60510e3",
x"d71ff0ef",
x"f59ff06f",
x"07500793",
x"02f41663",
x"ffe01537",
x"dd050513",
x"fccff0ef",
x"ffe005b7",
x"ffe00537",
x"15058593",
x"11850513",
x"fecff0ef",
x"0c050663",
x"00100073",
x"06500793",
x"00f41663",
x"d31ff0ef",
x"f25ff06f",
x"07800793",
x"fef404e3",
x"06800793",
x"00f41863",
x"ffe01537",
x"df050513",
x"f05ff06f",
x"06900793",
x"08f41663",
x"ffe01537",
x"e8050513",
x"f70ff0ef",
x"f1302573",
x"8c1ff0ef",
x"ffe01537",
x"e8850513",
x"f5cff0ef",
x"fffe0437",
x"00042503",
x"8a9ff0ef",
x"ffe01537",
x"e9050513",
x"f44ff0ef",
x"30102573",
x"895ff0ef",
x"ffe01537",
x"e9850513",
x"f30ff0ef",
x"fc002573",
x"881ff0ef",
x"ffe01537",
x"ea050513",
x"f1cff0ef",
x"00842503",
x"86dff0ef",
x"ffe01537",
x"ea850513",
x"f08ff0ef",
x"00442503",
x"859ff0ef",
x"ffe01537",
x"d2050513",
x"e75ff06f",
x"07300793",
x"02f40863",
x"06c00793",
x"e6f414e3",
x"ffe01537",
x"d8c50513",
x"ed8ff0ef",
x"ffe005b7",
x"ffe00537",
x"52c58593",
x"47050513",
x"ef8ff0ef",
x"e45ff06f",
x"800007b7",
x"0047a403",
x"00041863",
x"ffe01537",
x"eb050513",
x"e29ff06f",
x"929ff0ef",
x"00050863",
x"ffe01537",
x"c8450513",
x"e15ff06f",
x"ffe01537",
x"ec050513",
x"e88ff0ef",
x"00040513",
x"fd8ff0ef",
x"ffe01537",
x"ec850513",
x"e74ff0ef",
x"800004b7",
x"0004a503",
x"fc0ff0ef",
x"ffe01537",
x"edc50513",
x"e5cff0ef",
x"d8cff0ef",
x"07900793",
x"dcf51ae3",
x"ffe01537",
x"ee850513",
x"e44ff0ef",
x"01045413",
x"00140413",
x"004007b7",
x"00f4a023",
x"04041e63",
x"004007b7",
x"00f4a023",
x"0ff0000f",
x"0004a683",
x"00c68793",
x"00f4a023",
x"00000793",
x"80000737",
x"00472703",
x"06e7ee63",
x"b007c537",
x"0de50513",
x"00e12023",
x"00d4a023",
x"9b1ff0ef",
x"00012503",
x"9a9ff0ef",
x"fff44513",
x"9a1ff0ef",
x"ffe01537",
x"cc050513",
x"d59ff06f",
x"00600513",
x"00f12023",
x"ff8ff0ef",
x"f9cff0ef",
x"0d800513",
x"fd0ff0ef",
x"8bdff0ef",
x"facff0ef",
x"00012783",
x"fff40413",
x"00f12023",
x"ff8ff0ef",
x"00157513",
x"00012783",
x"fe0518e3",
x"00010737",
x"00e787b3",
x"f5dff06f",
x"00d12223",
x"0007a503",
x"00f12023",
x"00a40433",
x"939ff0ef",
x"00012783",
x"00412683",
x"00478793",
x"f5dff06f",
x"52524507",
x"445f524f",
x"43495645",
x"00000a45",
x"00000000",
x"52524507",
x"535f524f",
x"414e4749",
x"45525554",
x"0000000a",
x"52524507",
x"435f524f",
x"4b434548",
x"0a4d5553",
x"00000000",
x"000a4b4f",
x"5b1b070a",
x"31333b31",
x"5252456d",
x"455f524f",
x"50454358",
x"4e4f4954",
x"00000020",
x"6d305b1b",
x"0000000a",
x"65206f4e",
x"75636578",
x"6c626174",
x"42202e65",
x"20746f6f",
x"77796e61",
x"203f7961",
x"6e2f7928",
x"00000a29",
x"746f6f42",
x"20676e69",
x"6d6f7266",
x"00000020",
x"0a2e2e2e",
x"0000000a",
x"4e0a0a0a",
x"56524f45",
x"42203233",
x"6c746f6f",
x"6564616f",
x"75620a72",
x"3a646c69",
x"6e614a20",
x"20323220",
x"36323032",
x"00000a0a",
x"6f747541",
x"6f6f622d",
x"00000074",
x"206e6920",
x"202e7338",
x"73657250",
x"6e612073",
x"656b2079",
x"6f742079",
x"6f626120",
x"0a2e7472",
x"00000000",
x"726f6241",
x"2e646574",
x"00000a0a",
x"64616f4c",
x"20676e69",
x"6d6f7266",
x"49505320",
x"616c6620",
x"40206873",
x"30307830",
x"30303034",
x"2e2e3030",
x"0000202e",
x"65707954",
x"27682720",
x"726f6620",
x"6c656820",
x"000a2e70",
x"3a444d43",
x"0000203e",
x"69617741",
x"676e6974",
x"6f656e20",
x"32337672",
x"6578655f",
x"6e69622e",
x"202e2e2e",
x"00000000",
x"69617641",
x"6c62616c",
x"4d432065",
x"0a3a7344",
x"48203a68",
x"0a706c65",
x"53203a69",
x"65747379",
x"6e69206d",
x"720a6f66",
x"6552203a",
x"72617473",
x"3a750a74",
x"6c705520",
x"2064616f",
x"20616976",
x"54524155",
x"203a6c0a",
x"20495053",
x"73616c66",
x"202d2068",
x"64616f6c",
x"203a730a",
x"20495053",
x"73616c66",
x"202d2068",
x"676f7270",
x"0a6d6172",
x"53203a65",
x"74726174",
x"65786520",
x"61747563",
x"0a656c62",
x"45203a78",
x"0a746978",
x"00000000",
x"3a565748",
x"00002020",
x"4b4c430a",
x"0020203a",
x"53494d0a",
x"00203a41",
x"5349580a",
x"00203a41",
x"434f530a",
x"0020203a",
x"53494d0a",
x"00203a43",
x"65206f4e",
x"75636578",
x"6c626174",
x"000a2e65",
x"74697257",
x"00002065",
x"74796220",
x"74207365",
x"6c66206f",
x"20687361",
x"00000040",
x"7928203f",
x"0a296e2f",
x"00000000",
x"73616c46",
x"676e6968",
x"202e2e2e",
x"00000000",
x"33323130",
x"37363534",
x"62613938",
x"66656463",
others => (others => '0')
);

end neorv32_bootrom_image;
