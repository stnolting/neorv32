library ieee;
use ieee.std_logic_1164.all;

package neorv32_imem_image is

type rom_t is array (0 to 255) of std_ulogic_vector(31 downto 0);
constant image_size_c : natural := 772;
constant image_data_c : rom_t := (
x"f14020f3",
x"80002217",
x"ffb20213",
x"ff027113",
x"80000197",
x"7f018193",
x"000022b7",
x"80028293",
x"30029073",
x"00000317",
x"19030313",
x"30531073",
x"30401073",
x"00000397",
x"2d038393",
x"80000417",
x"fc440413",
x"80000497",
x"fbc48493",
x"80000517",
x"fb450513",
x"80000597",
x"fac58593",
x"00000613",
x"00000693",
x"00000713",
x"00000793",
x"00000813",
x"00000893",
x"00000913",
x"00000993",
x"00000a13",
x"00000a93",
x"00000b13",
x"00000b93",
x"00000c13",
x"00000c93",
x"00000d13",
x"00000d93",
x"00000e13",
x"00000e93",
x"00000f13",
x"00000f93",
x"04008263",
x"00000797",
x"01c78793",
x"30579073",
x"30445073",
x"30046073",
x"10500073",
x"ffdff06f",
x"00000797",
x"0e878793",
x"30579073",
x"fff44737",
x"00872103",
x"00c72603",
x"fff40737",
x"00072223",
x"05c0006f",
x"00838e63",
x"00945c63",
x"0003a783",
x"00f42023",
x"00438393",
x"00440413",
x"fedff06f",
x"00b55863",
x"00052023",
x"00450513",
x"ff5ff06f",
x"00000417",
x"1e840413",
x"00000497",
x"1e048493",
x"00945a63",
x"00042083",
x"000080e7",
x"00440413",
x"ff1ff06f",
x"00000617",
x"08c60613",
x"0ff0000f",
x"0000100f",
x"00000513",
x"00000593",
x"000600e7",
x"30047073",
x"30401073",
x"00000597",
x"05058593",
x"30559073",
x"34051073",
x"f1402473",
x"02041463",
x"00000417",
x"18840413",
x"00000497",
x"18048493",
x"00945a63",
x"00042083",
x"000080e7",
x"00440413",
x"ff1ff06f",
x"f1402473",
x"00041463",
x"00100073",
x"10500073",
x"ffdff06f",
x"10500073",
x"ffdff06f",
x"fffe07b7",
x"00050593",
x"0007a503",
x"0340006f",
x"ff010113",
x"00000513",
x"00812423",
x"00112623",
x"00000413",
x"064000ef",
x"0ff47513",
x"05c000ef",
x"0fa00513",
x"fcdff0ef",
x"00140413",
x"fedff06f",
x"ff010113",
x"00058613",
x"00000693",
x"00a55513",
x"00000593",
x"00112623",
x"060000ef",
x"01c59593",
x"00455513",
x"00a58533",
x"00050a63",
x"00001863",
x"fff50513",
x"00000013",
x"ff1ff06f",
x"00c12083",
x"01010113",
x"00008067",
x"fffc07b7",
x"00a7a223",
x"00008067",
x"00050613",
x"00000513",
x"0015f693",
x"00068463",
x"00c50533",
x"0015d593",
x"00161613",
x"fe0596e3",
x"00008067",
x"ff010113",
x"00068293",
x"00112623",
x"00050393",
x"00050693",
x"00060713",
x"00000793",
x"00000313",
x"00000813",
x"00d808b3",
x"00177e93",
x"00f30f33",
x"01f6de13",
x"00175713",
x"0108bfb3",
x"00179793",
x"000e8663",
x"00088813",
x"01ef8333",
x"00169693",
x"01c7e7b3",
x"fc0718e3",
x"00058863",
x"00060513",
x"f7dff0ef",
x"00650333",
x"00028a63",
x"00038513",
x"00028593",
x"f69ff0ef",
x"00650333",
x"00c12083",
x"00080513",
x"00030593",
x"01010113",
x"00008067",
others => (others => '0')
);

end neorv32_imem_image;
