-- #################################################################################################
-- # << NEORV32 - Custom Functions Subsystem (CFS) >>                                              #
-- # ********************************************************************************************* #
-- # Intended for tightly-coupled, application-specific custom co-processors. This module provides #
-- # 64x 32-bit memory-mapped interface registers, one interrupt request signal and custom IO      #
-- # conduits for processor-external or chip-external interface.                                   #
-- #                                                                                               #
-- # NOTE: This is just an example/illustration template. Modify/replace this file to implement    #
-- #       your own custom design logic.                                                           #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2022, Stephan Nolting. All rights reserved.                                     #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # The NEORV32 Processor - https://github.com/stnolting/neorv32              (c) Stephan Nolting #
-- #################################################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library neorv32;
use neorv32.neorv32_package.all;

entity neorv32_cfs is
  generic (
    BASE_ADDR : std_ulogic_vector(31 downto 0); -- module base address
    CFS_CONFIG   : std_ulogic_vector(31 downto 0); -- custom CFS configuration generic
    CFS_IN_SIZE  : natural; -- size of CFS input conduit in bits
    CFS_OUT_SIZE : natural  -- size of CFS output conduit in bits
  );
  port (
    -- host access --
    clk_i       : in  std_ulogic; -- global clock line
    rstn_i      : in  std_ulogic; -- global reset line, low-active, use as async
    priv_i      : in  std_ulogic; -- current CPU privilege mode
    addr_i      : in  std_ulogic_vector(31 downto 0); -- address
    rden_i      : in  std_ulogic; -- read enable
    wren_i      : in  std_ulogic; -- word write enable
    data_i      : in  std_ulogic_vector(31 downto 0); -- data in
    data_o      : out std_ulogic_vector(31 downto 0); -- data out
    ack_o       : out std_ulogic; -- transfer acknowledge
    err_o       : out std_ulogic; -- transfer error
    -- clock generator --
    clkgen_en_o : out std_ulogic; -- enable clock generator
    clkgen_i    : in  std_ulogic_vector(07 downto 0); -- "clock" inputs
    -- interrupt --
    irq_o       : out std_ulogic; -- interrupt request
    -- custom io (conduits) --
    cfs_in_i    : in  std_ulogic_vector(CFS_IN_SIZE-1 downto 0);  -- custom inputs
    cfs_out_o   : out std_ulogic_vector(CFS_OUT_SIZE-1 downto 0)  -- custom outputs
  );
end neorv32_cfs;

architecture neorv32_cfs_rtl of neorv32_cfs is

  -- IO space: module base address --
  -- WARNING: Do not modify the CFS base address or the CFS' occupied address
  -- space as this might cause access collisions with other processor modules.
  constant hi_abb_c : natural := index_size_f(io_size_c)-1; -- high address boundary bit
  constant lo_abb_c : natural := index_size_f(cfs_size_c); -- low address boundary bit

  -- interface configuration
  constant cfs_reg0_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(0 * 4, lo_abb_c));
  constant cfs_reg1_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(1 * 4, lo_abb_c));
  constant cfs_reg2_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(2 * 4, lo_abb_c));
  constant cfs_reg3_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(3 * 4, lo_abb_c));
  constant cfs_reg4_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(4 * 4, lo_abb_c));
  constant cfs_reg5_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(5 * 4, lo_abb_c));
  constant cfs_reg6_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(6 * 4, lo_abb_c));
  constant cfs_reg7_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(7 * 4, lo_abb_c));
  constant cfs_reg8_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(8 * 4, lo_abb_c));
  constant cfs_reg9_offset_c      : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(9 * 4, lo_abb_c));
  constant cfs_reg10_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(10 * 4, lo_abb_c));
  constant cfs_reg11_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(11 * 4, lo_abb_c));
  constant cfs_reg12_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(12 * 4, lo_abb_c));
  constant cfs_reg13_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(13 * 4, lo_abb_c));
  constant cfs_reg14_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(14 * 4, lo_abb_c));
  constant cfs_reg15_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(15 * 4, lo_abb_c));
  constant cfs_reg16_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(16 * 4, lo_abb_c));
  constant cfs_reg17_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(17 * 4, lo_abb_c));
  constant cfs_reg18_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(18 * 4, lo_abb_c));
  constant cfs_reg19_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(19 * 4, lo_abb_c));
  constant cfs_reg20_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(20 * 4, lo_abb_c));
  constant cfs_reg21_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(21 * 4, lo_abb_c));
  constant cfs_reg22_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(22 * 4, lo_abb_c));
  constant cfs_reg23_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(23 * 4, lo_abb_c));
  constant cfs_reg24_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(24 * 4, lo_abb_c));
  constant cfs_reg25_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(25 * 4, lo_abb_c));
  constant cfs_reg26_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(26 * 4, lo_abb_c));
  constant cfs_reg27_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(27 * 4, lo_abb_c));
  constant cfs_reg28_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(28 * 4, lo_abb_c));
  constant cfs_reg29_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(29 * 4, lo_abb_c));
  constant cfs_reg30_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(30 * 4, lo_abb_c));
  constant cfs_reg31_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(31 * 4, lo_abb_c));
  constant cfs_reg32_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(32 * 4, lo_abb_c));
  constant cfs_reg33_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(33 * 4, lo_abb_c));
  constant cfs_reg34_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(34 * 4, lo_abb_c));
  constant cfs_reg35_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(35 * 4, lo_abb_c));
  constant cfs_reg36_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(36 * 4, lo_abb_c));
  constant cfs_reg37_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(37 * 4, lo_abb_c));
  constant cfs_reg38_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(38 * 4, lo_abb_c));
  constant cfs_reg39_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(39 * 4, lo_abb_c));
  constant cfs_reg40_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(40 * 4, lo_abb_c));
  constant cfs_reg41_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(41 * 4, lo_abb_c));
  constant cfs_reg42_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(42 * 4, lo_abb_c));
  constant cfs_reg43_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(43 * 4, lo_abb_c));
  constant cfs_reg44_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(44 * 4, lo_abb_c));
  constant cfs_reg45_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(45 * 4, lo_abb_c));
  constant cfs_reg46_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(46 * 4, lo_abb_c));
  constant cfs_reg47_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(47 * 4, lo_abb_c));
  constant cfs_reg48_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(48 * 4, lo_abb_c));
  constant cfs_reg49_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(49 * 4, lo_abb_c));
  constant cfs_reg50_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(50 * 4, lo_abb_c));
  constant cfs_reg51_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(51 * 4, lo_abb_c));
  constant cfs_reg52_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(52 * 4, lo_abb_c));
  constant cfs_reg53_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(53 * 4, lo_abb_c));
  constant cfs_reg54_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(54 * 4, lo_abb_c));
  constant cfs_reg55_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(55 * 4, lo_abb_c));
  constant cfs_reg56_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(56 * 4, lo_abb_c));
  constant cfs_reg57_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(57 * 4, lo_abb_c));
  constant cfs_reg58_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(58 * 4, lo_abb_c));
  constant cfs_reg59_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(59 * 4, lo_abb_c));
  constant cfs_reg60_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(60 * 4, lo_abb_c));
  constant cfs_reg61_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(61 * 4, lo_abb_c));
  constant cfs_reg62_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(62 * 4, lo_abb_c));
  constant cfs_reg63_offset_c     : std_ulogic_vector(lo_abb_c-1 downto 0) := std_ulogic_vector(to_signed(63 * 4, lo_abb_c));

  -- access control --
  signal acc_en : std_ulogic; -- module access enable
  signal offset : std_ulogic_vector(lo_abb_c-1 downto 0); -- access address
  signal wren   : std_ulogic; -- word write enable
  signal rden   : std_ulogic; -- read enable

  -- default CFS interface registers --
  type cfs_regs_t is array (0 to 3) of std_ulogic_vector(31 downto 0); -- just implement 4 registers for this example
  signal cfs_reg_wr : cfs_regs_t; -- interface registers for WRITE accesses
  signal cfs_reg_rd : cfs_regs_t; -- interface registers for READ accesses

begin

  -- Access Control -------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- This logic is required to handle the CPU accesses - DO NOT MODIFY!
  acc_en <= '1' when (addr_i(hi_abb_c downto lo_abb_c) = BASE_ADDR(hi_abb_c downto lo_abb_c)) else '0';
  offset <= addr_i(lo_abb_c-1 downto 2) & "00"; -- word aligned
  wren   <= acc_en and wren_i; -- only full-word write accesses are supported
  rden   <= acc_en and rden_i; -- read accesses always return a full 32-bit word


  -- CFS Generics ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- In it's default version the CFS provides three configuration generics:
  -- > CFS_IN_SIZE  - configures the size (in bits) of the CFS input conduit cfs_in_i
  -- > CFS_OUT_SIZE - configures the size (in bits) of the CFS output conduit cfs_out_o
  -- > CFS_CONFIG   - is a blank 32-bit generic. It is intended as a "generic conduit" to propagate
  --                  custom configuration flags from the top entity down to this module.


  -- CFS IOs --------------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- By default, the CFS provides two IO signals (cfs_in_i and cfs_out_o) that are available at the processor's top entity.
  -- These are intended as "conduits" to propagate custom signals from this module and the processor top entity.

  cfs_out_o <= (others => '0'); -- not used for this minimal example


  -- Reset System ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- The CFS can be reset using the global rstn_i signal. This signal should be used as asynchronous reset and is active-low.
  -- Note that rstn_i can be asserted by a processor-external reset, the on-chip debugger and also by the watchdog.
  --
  -- Most default peripheral devices of the NEORV32 do NOT use a dedicated hardware reset at all. Instead, these units are
  -- reset by writing ZERO to a specific "control register" located right at the beginning of the device's address space
  -- (so this register is cleared at first). The crt0 start-up code writes ZERO to every single address in the processor's
  -- IO space - including the CFS. Make sure that this initial clearing does not cause any unintended CFS actions.


  -- Clock System ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- The processor top unit implements a clock generator providing 8 "derived clocks".
  -- Actually, these signals should not be used as direct clock signals, but as *clock enable* signals.
  -- clkgen_i is always synchronous to the main system clock (clk_i).
  --
  -- The following clock dividers are available:
  -- > clkgen_i(clk_div2_c)    -> MAIN_CLK/2
  -- > clkgen_i(clk_div4_c)    -> MAIN_CLK/4
  -- > clkgen_i(clk_div8_c)    -> MAIN_CLK/8
  -- > clkgen_i(clk_div64_c)   -> MAIN_CLK/64
  -- > clkgen_i(clk_div128_c)  -> MAIN_CLK/128
  -- > clkgen_i(clk_div1024_c) -> MAIN_CLK/1024
  -- > clkgen_i(clk_div2048_c) -> MAIN_CLK/2048
  -- > clkgen_i(clk_div4096_c) -> MAIN_CLK/4096
  --
  -- For instance, if you want to drive a clock process at MAIN_CLK/8 clock speed you can use the following construct:
  --
  --   if (rstn_i = '0') then -- async and low-active reset (if required at all)
  --   ...
  --   elsif rising_edge(clk_i) then -- always use the main clock for all clock processes
  --     if (clkgen_i(clk_div8_c) = '1') then -- the div8 "clock" is actually a clock enable
  --       ...
  --     end if;
  --   end if;
  --
  -- The clkgen_i input clocks are available when at least one IO/peripheral device (for example UART0) requires the clocks
  -- generated by the clock generator. The CFS can enable the clock generator by itself by setting the clkgen_en_o signal high.
  -- The CFS cannot ensure to deactivate the clock generator by setting the clkgen_en_o signal low as other peripherals might
  -- still keep the generator activated. Make sure to deactivate the CFS's clkgen_en_o if no clocks are required in here to
  -- reduce dynamic power consumption.

  clkgen_en_o <= '0'; -- not used for this minimal example


  -- Interrupt ------------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- The CFS features a single interrupt signal, which is connected to the CPU's "fast interrupt" channel 1 (FIRQ1).
  -- The interrupt is triggered by a one-cycle high-level. After triggering, the interrupt appears as "pending" in the CPU's
  -- mip CSR ready to trigger execution of the according interrupt handler. It is the task of the application to programmer
  -- to enable/clear the CFS interrupt using the CPU's mie and mip registers when required.

  irq_o <= '0'; -- not used for this minimal example


  -- Read/Write Access ----------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- Here we are reading/writing from/to the interface registers of the module and generate the CPU access handshake (bus response).
  --
  -- The CFS provides up to 64 memory-mapped 32-bit interface registers. For instance, these could be used to provide a
  -- <control register> for global control of the unit, a <data register> for reading/writing from/to a data FIFO, a
  -- <command register> for issuing commands and a <status register> for status information.
  --
  -- Following the interface protocol, each read or write access has to be acknowledged in the following cycle using the ack_o
  -- signal (or even later if the module needs additional time). If no ACK is generated at all, the bus access will time out
  -- and cause a bus access fault exception. The current CPU privilege level is available via the 'priv_i' signal (0 = user mode,
  -- 1 = machine mode), which can be used to constrain access to certain registers or features to privileged software only.
  --
  -- This module also provides an optional ERROR signal to indicate a faulty access operation (for example when accessing an
  -- unused, read-only or "locked" CFS register address). This signal may only be set when the module is actually accessed
  -- and is set INSTEAD of the ACK signal. Setting the ERR signal will raise a bus access exception with a "Device Error" qualifier
  -- that can be handled by the application software. Note that the current privilege level should not be exposed to software to
  -- maintain full virtualization. Hence, CFS-based "privilege escalation" should trigger a bus access exception (e.g. by setting 'err_o').

  err_o <= '0'; -- Tie to zero if not explicitly used.


  -- Host access example: Read and write access to the interface registers + bus transfer acknowledge. This example only
  -- implements four physical r/w register (the four lowest CFS registers). The remaining addresses of the CFS are not associated
  -- with any physical registers - any access to those is simply ignored but still acknowledged. Only full-word write accesses are
  -- supported (and acknowledged) by this example. Sub-word write access will not alter any CFS register state and will cause
  -- a "bus store access" exception (with a "Device Timeout" qualifier as not ACK is generated in that case).

  host_access: process(rstn_i, clk_i)
  begin
    if (rstn_i = '0') then
      cfs_reg_wr(0) <= (others => '0');
      cfs_reg_wr(1) <= (others => '0');
      cfs_reg_wr(2) <= (others => '0');
      cfs_reg_wr(3) <= (others => '0');
      --
      ack_o  <= '0';
      data_o <= (others => '0');
    elsif rising_edge(clk_i) then -- synchronous interface for read and write accesses
      -- transfer/access acknowledge --
      -- default: required for the CPU to check the CFS is answering a bus read OR write request;
      -- all read and write accesses (to any cfs_reg, even if there is no according physical register implemented) will succeed.
      ack_o <= rden or wren;

      -- write access --
      if (wren = '1') then -- full-word write access, high for one cycle if there is an actual write access
        if (offset = cfs_reg0_offset_c) then -- make sure to use the internal "offset" signal for the read/write interface
          cfs_reg_wr(0) <= data_i; -- some physical register, for example: control register
        end if;
        if (offset = cfs_reg1_offset_c) then
          cfs_reg_wr(1) <= data_i; -- some physical register, for example: data in/out fifo
        end if;
        if (offset = cfs_reg2_offset_c) then
          cfs_reg_wr(2) <= data_i; -- some physical register, for example: command fifo
        end if;
        if (offset = cfs_reg3_offset_c) then
          cfs_reg_wr(3) <= data_i; -- some physical register, for example: status register
        end if;
      end if;

      -- read access --
      data_o <= (others => '0'); -- the output HAS TO BE ZERO if there is no actual read access
      if (rden = '1') then -- the read access is always 32-bit wide, high for one cycle if there is an actual read access
        case offset is -- make sure to use the internal 'offset' signal for the read/write interface
          when cfs_reg0_offset_c => data_o <= cfs_reg_rd(0);
          when cfs_reg1_offset_c => data_o <= cfs_reg_rd(1);
          when cfs_reg2_offset_c => data_o <= cfs_reg_rd(2);
          when cfs_reg3_offset_c => data_o <= cfs_reg_rd(3);
          when others          => data_o <= (others => '0'); -- the remaining registers are not implemented and will read as zero
        end case;
      end if;
    end if;
  end process host_access;


  -- CFS Function Core ----------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------

  -- This is where the actual functionality can be implemented.
  -- The logic below is just a very simple example that transforms data
  -- from an input register into data in an output register.

  cfs_reg_rd(0) <= bin_to_gray_f(cfs_reg_wr(0)); -- convert binary to gray code
  cfs_reg_rd(1) <= gray_to_bin_f(cfs_reg_wr(1)); -- convert gray to binary code
  cfs_reg_rd(2) <= bit_rev_f(cfs_reg_wr(2)); -- bit reversal
  cfs_reg_rd(3) <= bswap32_f(cfs_reg_wr(3)); -- byte swap (endianness conversion)


end neorv32_cfs_rtl;
