-- #################################################################################################
-- # << NEORV32 - Default Testbench >>                                                             #
-- # ********************************************************************************************* #
-- # This testbench provides a virtual UART receiver connected to the processor's uart_txd_o       #
-- # signal. The received chars are shown in the simulator console and also written to a file      #
-- # ("neorv32.testbench_uart.out"). Futhermore, this testbench provides a simple RAM connected    #
-- # to the external Wishbone bus. The testbench configures the processor with all optional        #
-- # elements enabled by default.                                                                  #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2020, Stephan Nolting. All rights reserved.                                     #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # The NEORV32 Processor - https://github.com/stnolting/neorv32              (c) Stephan Nolting #
-- #################################################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library neorv32;
use neorv32.neorv32_package.all;
use neorv32.neorv32_application_image.all; -- this file is generated by the image generator
use std.textio.all;

entity neorv32_tb is
end neorv32_tb;

architecture neorv32_tb_rtl of neorv32_tb is

  -- User Configuration ---------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant t_clock_c          : time := 10 ns; -- main clock period
  constant f_clock_c          : real := 100000000.0; -- main clock in Hz
  constant f_clock_nat_c      : natural := 100000000; -- main clock in Hz
  constant baud_rate_c        : real := 19200.0; -- standard UART baudrate
  --
  constant wb_mem_base_addr_c : std_ulogic_vector(31 downto 0) := x"F0000000"; -- wishbone memory base address
  constant wb_mem_size_c      : natural := 256; -- wishbone memory size in bytes
  constant wb_mem_latency_c   : natural := 8; -- latency in clock cycles (min 1)
  -- -------------------------------------------------------------------------------------------

  -- text.io --
  file file_uart_tx_out : text open write_mode is "neorv32.testbench_uart.out";

  -- internal configuration --
  constant baud_val_c : real    := f_clock_c / baud_rate_c;
  constant f_clk_c    : natural := natural(f_clock_c);

  -- generators --
  signal clk_gen, rst_gen : std_ulogic := '0';

  -- simulation uart receiver --
  signal uart_txd         : std_ulogic;
  signal uart_rx_sync     : std_ulogic_vector(04 downto 0) := (others => '1');
  signal uart_rx_busy     : std_ulogic := '0';
  signal uart_rx_sreg     : std_ulogic_vector(08 downto 0) := (others => '0');
  signal uart_rx_baud_cnt : real;
  signal uart_rx_bitcnt   : natural;

  -- gpio --
  signal gpio : std_ulogic_vector(31 downto 0);

  -- twi --
  signal twi_scl, twi_sda : std_logic;

  -- spi --
  signal spi_data : std_logic;

  -- Wishbone bus --
  type wishbone_t is record
    addr  : std_ulogic_vector(31 downto 0); -- address
    wdata : std_ulogic_vector(31 downto 0); -- master write data
    rdata : std_ulogic_vector(31 downto 0); -- master read data
    we    : std_ulogic; -- write enable
    sel   : std_ulogic_vector(03 downto 0); -- byte enable
    stb   : std_ulogic; -- strobe
    cyc   : std_ulogic; -- valid cycle
    ack   : std_ulogic; -- transfer acknowledge
    err   : std_ulogic; -- transfer error
    tag   : std_ulogic_vector(2 downto 0); -- tag
  end record;
  signal wb_cpu : wishbone_t;

  -- Wishbone memory --
  type wb_mem_ram_t is array (0 to wb_mem_size_c/4-1) of std_ulogic_vector(31 downto 0);
  type wb_mem_read_latency_t is array (0 to wb_mem_latency_c-1) of std_ulogic_vector(31 downto 0);

  -- init function --
  -- impure function: returns NOT the same result every time it is evaluated with the same arguments since the source file might have changed
  impure function init_wbmem(init : application_init_image_t) return wb_mem_ram_t is
    variable mem_v : wb_mem_ram_t;
  begin
    mem_v := (others => (others => '0'));
    for i in 0 to init'length-1 loop -- init only in range of source data array
        mem_v(i) := init(i);
    end loop; -- i
    return mem_v;
  end function init_wbmem;

  -- ---------------------------------------------- --
  -- How to simulate a boot from an external memory --
  -- ---------------------------------------------- --
  -- The simulated Wishbone memory can be initialized with the compiled application init.
  -- 1. Uncomment the init_wbmem function below; this will initialize the simulated wishbone memory with the neorv32_application_image.vhd image
  -- 2. Increase the wb_mem_size_c constant above to (at least) the size of the application image (like 16kB -> 16*1024)
  -- 3. Disable the processor-internal IMEM in the processor instantiation below (MEM_INT_IMEM_USE => false)
  -- 4. Set the Wishbone memory base address wb_mem_base_addr_c (above) to zero (constant wb_mem_base_addr_c : std_ulogic_vector(31 downto 0) := x"00000000";)
  -- 5. Simulate!

  signal wb_ram : wb_mem_ram_t;-- := init_wbmem(application_init_image); -- uncomment if you want to init the WB ram with app image

  type wb_mem_t is record
    rdata  : wb_mem_read_latency_t;
    acc_en : std_ulogic;
    ack    : std_ulogic_vector(wb_mem_latency_c-1 downto 0);
    rb_en  : std_ulogic_vector(wb_mem_latency_c-1 downto 0);
  end record;
  signal wb_mem : wb_mem_t;

begin

  -- Clock/Reset Generator ------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  clk_gen <= not clk_gen after (t_clock_c/2);
  rst_gen <= '0', '1' after 60*(t_clock_c/2);


  -- CPU Core -------------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  neorv32_top_inst: neorv32_top
  generic map (
    -- General --
    CLOCK_FREQUENCY              => f_clock_nat_c, -- clock frequency of clk_i in Hz
    BOOTLOADER_USE               => false,         -- implement processor-internal bootloader?
    USER_CODE                    => x"12345678",   -- custom user code
    -- RISC-V CPU Extensions --
    CPU_EXTENSION_RISCV_C        => true,          -- implement compressed extension?
    CPU_EXTENSION_RISCV_E        => false,         -- implement embedded RF extension?
    CPU_EXTENSION_RISCV_M        => true,          -- implement muld/div extension?
    CPU_EXTENSION_RISCV_U        => true,          -- implement user mode extension?
    CPU_EXTENSION_RISCV_Zicsr    => true,          -- implement CSR system?
    CPU_EXTENSION_RISCV_Zifencei => true,          -- implement instruction stream sync.?
    -- Extension Options --
    FAST_MUL_EN                  => false,         -- use DSPs for M extension's multiplier
    FAST_SHIFT_EN                => false,         -- use barrel shifter for shift operations
    -- Physical Memory Protection (PMP) --
    PMP_USE                      => true,          -- implement PMP?
    PMP_NUM_REGIONS              => 4,             -- number of regions (max 16)
    PMP_GRANULARITY              => 14,            -- minimal region granularity (1=8B, 2=16B, 3=32B, ...) default is 64k
    -- Internal Instruction memory --
    MEM_INT_IMEM_USE             => true,          -- implement processor-internal instruction memory
    MEM_INT_IMEM_SIZE            => 16*1024,       -- size of processor-internal instruction memory in bytes
    MEM_INT_IMEM_ROM             => false,         -- implement processor-internal instruction memory as ROM
    -- Internal Data memory --
    MEM_INT_DMEM_USE             => true,          -- implement processor-internal data memory
    MEM_INT_DMEM_SIZE            => 8*1024,        -- size of processor-internal data memory in bytes
    -- External memory interface --
    MEM_EXT_USE                  => true,          -- implement external memory bus interface?
    -- Processor peripherals --
    IO_GPIO_USE                  => true,          -- implement general purpose input/output port unit (GPIO)?
    IO_MTIME_USE                 => true,          -- implement machine system timer (MTIME)?
    IO_UART_USE                  => true,          -- implement universal asynchronous receiver/transmitter (UART)?
    IO_SPI_USE                   => true,          -- implement serial peripheral interface (SPI)?
    IO_TWI_USE                   => true,          -- implement two-wire interface (TWI)?
    IO_PWM_USE                   => true,          -- implement pulse-width modulation unit (PWM)?
    IO_WDT_USE                   => true,          -- implement watch dog timer (WDT)?
    IO_TRNG_USE                  => false,         -- DEFAULT TRNG CONFIG CANNOT BE SIMULATED!
    IO_CFU0_USE                  => true,          -- implement custom functions unit 0 (CFU0)?
    IO_CFU1_USE                  => true           -- implement custom functions unit 1 (CFU1)?
  )
  port map (
    -- Global control --
    clk_i       => clk_gen,         -- global clock, rising edge
    rstn_i      => rst_gen,         -- global reset, low-active, async
    -- Wishbone bus interface --
    wb_tag_o    => wb_cpu.tag,      -- tag
    wb_adr_o    => wb_cpu.addr,     -- address
    wb_dat_i    => wb_cpu.rdata,    -- read data
    wb_dat_o    => wb_cpu.wdata,    -- write data
    wb_we_o     => wb_cpu.we,       -- read/write
    wb_sel_o    => wb_cpu.sel,      -- byte enable
    wb_stb_o    => wb_cpu.stb,      -- strobe
    wb_cyc_o    => wb_cpu.cyc,      -- valid cycle
    wb_ack_i    => wb_cpu.ack,      -- transfer acknowledge
    wb_err_i    => wb_cpu.err,      -- transfer error
    -- Advanced memory control signals --
    fence_o     => open,            -- indicates an executed FENCE operation
    fencei_o    => open,            -- indicates an executed FENCEI operation
    -- GPIO --
    gpio_o      => gpio,            -- parallel output
    gpio_i      => gpio,            -- parallel input
    -- UART --
    uart_txd_o  => uart_txd,        -- UART send data
    uart_rxd_i  => uart_txd,        -- UART receive data
    -- SPI --
    spi_sck_o   => open,            -- SPI serial clock
    spi_sdo_o   => spi_data,        -- controller data out, peripheral data in
    spi_sdi_i   => spi_data,        -- controller data in, peripheral data out
    spi_csn_o   => open,            -- SPI CS
    -- TWI --
    twi_sda_io  => twi_sda,         -- twi serial data line
    twi_scl_io  => twi_scl,         -- twi serial clock line
    -- PWM --
    pwm_o       => open,            -- pwm channels
    -- Interrupts --
    mtime_irq_i => '0',             -- machine software interrupt, available if IO_MTIME_USE = false
    msw_irq_i   => '0',             -- machine software interrupt
    mext_irq_i  => '0'              -- machine external interrupt
  );

  -- TWI termination (pull-ups) --
  twi_scl <= 'H';
  twi_sda <= 'H';


  -- Console UART Receiver ------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  uart_rx_console: process(clk_gen)
    variable i : integer;
    variable l : line;
  begin
    -- "UART" --
    if rising_edge(clk_gen) then
      -- synchronizer --
      uart_rx_sync <= uart_rx_sync(3 downto 0) & uart_txd;
      -- arbiter --
      if (uart_rx_busy = '0') then -- idle
        uart_rx_busy     <= '0';
        uart_rx_baud_cnt <= round(0.5 * baud_val_c);
        uart_rx_bitcnt   <= 9;
        if (uart_rx_sync(4 downto 1) = "1100") then -- start bit? (falling edge)
          uart_rx_busy <= '1';
        end if;
      else
        if (uart_rx_baud_cnt = 0.0) then
          if (uart_rx_bitcnt = 1) then
            uart_rx_baud_cnt <= round(0.5 * baud_val_c);
          else
            uart_rx_baud_cnt <= round(baud_val_c);
          end if;
          if (uart_rx_bitcnt = 0) then
            uart_rx_busy <= '0'; -- done
            i := to_integer(unsigned(uart_rx_sreg(8 downto 1)));

            if (i < 32) or (i > 32+95) then -- printable char?
              report "NEORV32_TB_UART.TX: (" & integer'image(i) & ")"; -- print code
            else
              report "NEORV32_TB_UART.TX: " & character'val(i); -- print ASCII
            end if;

            if (i = 10) then -- Linux line break
              writeline(file_uart_tx_out, l);
            elsif (i /= 13) then -- Remove additional carriage return
              write(l, character'val(i));
            end if;
          else
            uart_rx_sreg   <= uart_rx_sync(4) & uart_rx_sreg(8 downto 1);
            uart_rx_bitcnt <= uart_rx_bitcnt - 1;
          end if;
        else
          uart_rx_baud_cnt <= uart_rx_baud_cnt - 1.0;
        end if;
      end if;
    end if;
  end process uart_rx_console;


  -- Wishbone Memory (simulated external memory) --------------------------------------------
  -- -------------------------------------------------------------------------------------------
  wb_mem_ram_access: process(clk_gen)
  begin
    if rising_edge(clk_gen) then
      -- control --
      wb_mem.rb_en(0) <= wb_cpu.cyc and wb_cpu.stb and wb_mem.acc_en and (not wb_cpu.we); -- read-back control
      wb_mem.ack(0)   <= wb_cpu.cyc and wb_cpu.stb and wb_mem.acc_en; -- wishbone acknowledge
      -- write access --
      if ((wb_cpu.cyc and wb_cpu.stb and wb_mem.acc_en and wb_cpu.we) = '1') then -- valid write access
        for i in 0 to 3 loop
          if (wb_cpu.sel(i) = '1') then
            wb_ram(to_integer(unsigned(wb_cpu.addr(index_size_f(wb_mem_size_c/4)+1 downto 2))))(7+i*8 downto 0+i*8) <= wb_cpu.wdata(7+i*8 downto 0+i*8);
          end if;
        end loop; -- i
      end if;
      -- read access --
      wb_mem.rdata(0) <= wb_ram(to_integer(unsigned(wb_cpu.addr(index_size_f(wb_mem_size_c/4)+1 downto 2)))); -- word aligned
      -- virtual read and ack latency --
      if (wb_mem_latency_c > 1) then
        for i in 1 to wb_mem_latency_c-1 loop
          wb_mem.rdata(i) <= wb_mem.rdata(i-1);
          wb_mem.rb_en(i) <= wb_mem.rb_en(i-1) and wb_cpu.cyc;
          wb_mem.ack(i)   <= wb_mem.ack(i-1) and wb_cpu.cyc;
        end loop;
      end if;
    end if;
  end process wb_mem_ram_access;

  -- wishbone memory access? --
  wb_mem.acc_en <= '1' when (wb_cpu.addr >= wb_mem_base_addr_c) and (wb_cpu.addr < std_ulogic_vector(unsigned(wb_mem_base_addr_c) + wb_mem_size_c)) else '0';

  -- output to cpu --
  wb_cpu.rdata <= wb_mem.rdata(wb_mem_latency_c-1) when (wb_mem.rb_en(wb_mem_latency_c-1) = '1') else (others=> '0'); -- data output gate
  wb_cpu.ack   <= wb_mem.ack(wb_mem_latency_c-1);
  wb_cpu.err   <= '0';


end neorv32_tb_rtl;
