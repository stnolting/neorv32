-- #################################################################################################
-- # << NEORV32 - Example setup including the bootloader, for the TinyFPGA-BX (c) Board >>                #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2021, Stephan Nolting. All rights reserved.                                     #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # The NEORV32 Processor - https://github.com/stnolting/neorv32              (c) Stephan Nolting #
-- #################################################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library iCE40;
use iCE40.components.all; -- for device primitives and macros

entity neorv32_TinyFPGA_BX_BoardTop_MinimalBoot is
  port (
    -- 16 MHz Clock input
    TinyFPGABX_CLK   : in std_logic;
    -- LED outputs
    TinyFPGABX_LED   : out std_logic;
    -- USB Pins (which should be statically driven if not being used)
    TinyFPGABX_USBP  : out std_logic;
    TinyFPGABX_USBN  : out std_logic;
    TinyFPGABX_USBPU : out std_logic
  );
end entity;

architecture neorv32_TinyFPGA_BX_BoardTop_MinimalBoot_rtl of neorv32_TinyFPGA_BX_BoardTop_MinimalBoot is

  -- configuration --
  constant f_clock_c : natural := 20000000; -- PLL output clock frequency in Hz

  -- Globals
  signal pll_rstn : std_logic;
  signal pll_clk  : std_logic;

  -- internal IO connection --
  signal con_gpio_o : std_ulogic_vector(3 downto 0);

begin

  -- Assign USB pins to "0" so as to disconnect TinyFPGA-BX from
  -- the host system.  Otherwise it would try to talk to
  -- us over USB, which wouldn't work since we have no stack.
  TinyFPGABX_USBP  <= '0';
  TinyFPGABX_USBN  <= '0';
  TinyFPGABX_USBPU <= '0';


  -- System PLL -----------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- Settings generated by icepll -i 16 -o 20:
  -- F_PLLIN:      16.000 MHz (given)
  -- F_PLLOUT:     20.000 MHz (requested)
  -- F_PLLOUT:     20.000 MHz (achieved)
  -- FEEDBACK:     SIMPLE
  -- F_PFD:        16.000 MHz
  -- F_VCO:        640.000 MHz
  -- DIVR:         0 (4'b0000)
  -- DIVF:        39 (7'b0100111)
  -- DIVQ:         5 (3'b101)
  -- FILTER_RANGE: 1 (3'b001)
  Pll_inst : SB_PLL40_CORE
  generic map (
    FEEDBACK_PATH => "SIMPLE",
    DIVR          =>  x"0",
    DIVF          => 7x"27",
    DIVQ          => 3x"5",
    FILTER_RANGE  => 3x"1"
  )
  port map (
    REFERENCECLK    => TinyFPGABX_CLK,
    PLLOUTCORE      => open,
    PLLOUTGLOBAL    => pll_clk,
    EXTFEEDBACK     => '0',
    DYNAMICDELAY    => x"00",
    LOCK            => pll_rstn,
    BYPASS          => '0',
    RESETB          => '1',
    LATCHINPUTVALUE => '0',
    SDO             => open,
    SDI             => '0',
    SCLK            => '0'
  );

  -- The core of the problem ----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------

  neorv32_inst: entity work.neorv32_ProcessorTop_MinimalBoot
  generic map (
    CLOCK_FREQUENCY   => f_clock_c,  -- clock frequency of clk_i in Hz
    INT_BOOTLOADER_EN => true,
    MEM_INT_IMEM_EN   => false,
    MEM_INT_IMEM_SIZE => 8*1024,
    MEM_INT_DMEM_EN   => true,
    MEM_INT_DMEM_SIZE => 4*1024
  )
  port map (
    -- Global control --
    clk_i      => std_ulogic(pll_clk),
    rstn_i     => std_ulogic(pll_rstn),

    -- GPIO --
    gpio_o     => con_gpio_o,

    -- primary UART --
    uart_txd_o => open, -- UART0 send data
    uart_rxd_i => '0',  -- UART0 receive data
    uart_rts_o => open, -- hw flow control: UART0.RX ready to receive ("RTR"), low-active, optional
    uart_cts_i => '0',  -- hw flow control: UART0.TX allowed to transmit, low-active, optional

    -- PWM --
    pwm_o      => open
  );

  TinyFPGABX_LED <= con_gpio_o(0);

end architecture;
