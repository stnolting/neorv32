-- ================================================================================ --
-- NEORV32 SoC - Processor-internal bootloader ROM (BOOTROM)                        --
-- -------------------------------------------------------------------------------- --
-- The NEORV32 RISC-V Processor - https://github.com/stnolting/neorv32              --
-- Copyright (c) NEORV32 contributors.                                              --
-- Copyright (c) 2020 - 2024 Stephan Nolting. All rights reserved.                  --
-- Licensed under the BSD-3-Clause license, see LICENSE for details.                --
-- SPDX-License-Identifier: BSD-3-Clause                                            --
-- ================================================================================ --

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library neorv32;
use neorv32.neorv32_package.all;
use neorv32.neorv32_bootloader_image.all; -- this file is generated by the image generator

entity neorv32_boot_rom is
  port (
    clk_i     : in  std_ulogic; -- global clock line
    rstn_i    : in  std_ulogic; -- async reset, low-active
    bus_req_i : in  bus_req_t;  -- bus request
    bus_rsp_o : out bus_rsp_t   -- bus response
  );
end neorv32_boot_rom;

architecture neorv32_boot_rom_rtl of neorv32_boot_rom is

  -- determine physical ROM size in bytes (expand to next power of two) --
  constant boot_rom_size_index_c : natural := index_size_f((bootloader_init_size_c)); -- address with (bytes)
  constant boot_rom_size_c       : natural range 0 to iodev_size_c := (2**boot_rom_size_index_c); -- physical size in bytes

  -- ROM initialized with executable code --
  constant mem_rom_c : mem32_t(0 to boot_rom_size_c/4-1) := mem32_init_f(bootloader_init_image_c, boot_rom_size_c/4);

  -- local signals --
  signal rden  : std_ulogic;
  signal rdata : std_ulogic_vector(31 downto 0);

begin

  -- Memory Access --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  mem_access: process(clk_i)
  begin
    if rising_edge(clk_i) then -- no reset to infer block RAM
      rdata <= mem_rom_c(to_integer(unsigned(bus_req_i.addr(boot_rom_size_index_c+1 downto 2))));
    end if;
  end process mem_access;


  -- Bus Feedback ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  bus_feedback: process(rstn_i, clk_i)
  begin
    if (rstn_i = '0') then
      rden <= '0';
    elsif rising_edge(clk_i) then
      rden <= bus_req_i.stb and (not bus_req_i.rw); -- read-only
    end if;
  end process bus_feedback;

  bus_rsp_o.data <= rdata when (rden = '1') else (others => '0'); -- output gate
  bus_rsp_o.ack  <= rden;
  bus_rsp_o.err  <= '0'; -- no access error possible


end neorv32_boot_rom_rtl;
